// master.v

// Generated using ACDS version 13.1 162 at 2021.07.22.16:40:43

`timescale 1 ps / 1 ps
module master (
		input  wire        clk_50,                                                    //                               clk_50_clk_in.clk
		input  wire        reset_n,                                                   //                         clk_50_clk_in_reset.reset_n
		output wire [7:0]  pio_led_external_connection_export,                        //                 pio_led_external_connection.export
		output wire        commands_parameters_qsys_0_conduit_comm_par_start,         // commands_parameters_qsys_0_conduit_comm_par.start
		output wire        commands_parameters_qsys_0_conduit_comm_par_start_N,       //                                            .start_N
		output wire        commands_parameters_qsys_0_conduit_comm_par_auto,          //                                            .auto
		output wire        commands_parameters_qsys_0_conduit_comm_par_stop,          //                                            .stop
		input  wire [31:0] commands_parameters_qsys_0_conduit_comm_par_fi_phm,        //                                            .fi_phm
		input  wire [31:0] commands_parameters_qsys_0_conduit_comm_par_detuning,      //                                            .detuning
		input  wire        commands_parameters_qsys_0_conduit_comm_par_syncpulse,     //                                            .syncpulse
		input  wire        commands_parameters_qsys_0_conduit_comm_par_TURN_ON_RF,    //                                            .TURN_ON_RF
		output wire [31:0] commands_parameters_qsys_0_conduit_comm_par_d_fi_gate2,    //                                            .d_fi_gate2
		output wire [31:0] commands_parameters_qsys_0_conduit_comm_par_d_i_gate2,     //                                            .d_i_gate2
		output wire [31:0] commands_parameters_qsys_0_conduit_comm_par_dx2,           //                                            .dx2
		output wire [31:0] commands_parameters_qsys_0_conduit_comm_par_dx1,           //                                            .dx1
		output wire [31:0] commands_parameters_qsys_0_conduit_comm_par_DZ_TP,         //                                            .DZ_TP
		output wire [31:0] commands_parameters_qsys_0_conduit_comm_par_DZ_TX,         //                                            .DZ_TX
		output wire [31:0] commands_parameters_qsys_0_conduit_comm_par_PULSE_NUMBER,  //                                            .PULSE_NUMBER
		output wire [31:0] commands_parameters_qsys_0_conduit_comm_par_DZ_TR,         //                                            .DZ_TR
		output wire [31:0] commands_parameters_qsys_0_conduit_comm_par_period_MANUAL, //                                            .period_MANUAL
		output wire [31:0] commands_parameters_qsys_0_conduit_comm_par_L,             //                                            .L
		output wire [31:0] commands_parameters_qsys_0_conduit_comm_par_F2,            //                                            .F2
		output wire [31:0] commands_parameters_qsys_0_conduit_comm_par_F1,            //                                            .F1
		output wire        commands_parameters_qsys_0_conduit_comm_par_count_MANUAL,  //                                            .count_MANUAL
		output wire        commands_parameters_qsys_0_conduit_comm_par_dir_MANUAL,    //                                            .dir_MANUAL
		output wire        commands_parameters_qsys_0_conduit_comm_par_tp,            //                                            .tp
		output wire        commands_parameters_qsys_0_conduit_comm_par_tx,            //                                            .tx
		output wire        commands_parameters_qsys_0_conduit_comm_par_tr,            //                                            .tr
		input  wire [15:0] commands_parameters_qsys_0_s0_address,                     //               commands_parameters_qsys_0_s0.address
		input  wire [31:0] commands_parameters_qsys_0_s0_writedata,                   //                                            .writedata
		output wire [31:0] commands_parameters_qsys_0_s0_readdata,                    //                                            .readdata
		input  wire        commands_parameters_qsys_0_s0_write,                       //                                            .write
		input  wire        commands_parameters_qsys_0_s0_read,                        //                                            .read
		output wire [31:0] pulse_qsys_conduit_drv_pulse,                              //                          pulse_qsys_conduit.drv_pulse
		input  wire        pulse_qsys_conduit_drv_dir,                                //                                            .drv_dir
		input  wire        pulse_qsys_conduit_enable,                                 //                                            .enable
		input  wire        pulse_qsys_conduit_counter_en,                             //                                            .counter_en
		input  wire [31:0] pulse_qsys_conduit_drv_period,                             //                                            .drv_period
		input  wire [31:0] pulse_qsys_conduit_PULSE_NUMBER,                           //                                            .PULSE_NUMBER
		output wire [31:0] mux_qsys_conduit_drv_period,                               //                            mux_qsys_conduit.drv_period
		output wire        mux_qsys_conduit_drv_dir,                                  //                                            .drv_dir
		output wire        mux_qsys_conduit_enable,                                   //                                            .enable
		output wire        mux_qsys_conduit_counter_en,                               //                                            .counter_en
		input  wire [31:0] mux_qsys_conduit_period_TR,                                //                                            .period_TR
		input  wire [31:0] mux_qsys_conduit_period_TX,                                //                                            .period_TX
		input  wire [31:0] mux_qsys_conduit_period_TP,                                //                                            .period_TP
		input  wire [31:0] mux_qsys_conduit_detuning,                                 //                                            .detuning
		input  wire [31:0] mux_qsys_conduit_fi_phm,                                   //                                            .fi_phm
		input  wire        mux_qsys_conduit_tr,                                       //                                            .tr
		input  wire        mux_qsys_conduit_tx,                                       //                                            .tx
		input  wire        mux_qsys_conduit_tp,                                       //                                            .tp
		input  wire        mux_qsys_conduit_dir_TX,                                   //                                            .dir_TX
		input  wire        mux_qsys_conduit_dir_TR,                                   //                                            .dir_TR
		input  wire        mux_qsys_conduit_dir_TP,                                   //                                            .dir_TP
		input  wire        mux_qsys_conduit_drv_en_TR,                                //                                            .drv_en_TR
		input  wire        mux_qsys_conduit_drv_en_TX,                                //                                            .drv_en_TX
		input  wire        mux_qsys_conduit_drv_en_TP,                                //                                            .drv_en_TP
		input  wire        mux_qsys_conduit_counter_en_TR,                            //                                            .counter_en_TR
		input  wire        mux_qsys_conduit_syncpulse,                                //                                            .syncpulse
		input  wire [15:0] tp_qsys_conduit_k_TP,                                      //                             tp_qsys_conduit.k_TP
		input  wire [15:0] tp_qsys_conduit_d_fi_gate2,                                //                                            .d_fi_gate2
		input  wire [15:0] tp_qsys_conduit_L,                                         //                                            .L
		input  wire [15:0] tp_qsys_conduit_DZ_TP,                                     //                                            .DZ_TP
		input  wire [15:0] tp_qsys_conduit_F2,                                        //                                            .F2
		input  wire [15:0] tp_qsys_conduit_F1,                                        //                                            .F1
		input  wire [15:0] tp_qsys_conduit_detuning,                                  //                                            .detuning
		input  wire [15:0] tp_qsys_conduit_fi_set,                                    //                                            .fi_set
		input  wire [15:0] tp_qsys_conduit_fi_phm,                                    //                                            .fi_phm
		input  wire        tp_qsys_conduit_tp_mode,                                   //                                            .tp_mode
		input  wire        tp_qsys_conduit_data_valid_TP,                             //                                            .data_valid_TP
		output wire [31:0] tp_qsys_conduit_period_TP,                                 //                                            .period_TP
		output wire        tp_qsys_conduit_dir_TP,                                    //                                            .dir_TP
		output wire        tp_qsys_conduit_drv_en_TP,                                 //                                            .drv_en_TP
		input  wire        tx_qsys_conduit_syncpulse,                                 //                             tx_qsys_conduit.syncpulse
		input  wire [19:0] tx_qsys_conduit_k_TX,                                      //                                            .k_TX
		input  wire [15:0] tx_qsys_conduit_d_i_gate2,                                 //                                            .d_i_gate2
		input  wire [15:0] tx_qsys_conduit_DZ_TX,                                     //                                            .DZ_TX
		input  wire [15:0] tx_qsys_conduit_L,                                         //                                            .L
		input  wire [15:0] tx_qsys_conduit_F2,                                        //                                            .F2
		input  wire [15:0] tx_qsys_conduit_F1,                                        //                                            .F1
		input  wire [15:0] tx_qsys_conduit_i_fid_TX,                                  //                                            .i_fid_TX
		input  wire [15:0] tx_qsys_conduit_i_set,                                     //                                            .i_set
		input  wire        tx_qsys_conduit_tx_mode,                                   //                                            .tx_mode
		input  wire [15:0] tx_qsys_conduit_i_fid,                                     //                                            .i_fid
		input  wire        tx_qsys_conduit_data_valid_TX,                             //                                            .data_valid_TX
		output wire [31:0] tx_qsys_conduit_period_TX,                                 //                                            .period_TX
		output wire        tx_qsys_conduit_dir_TX,                                    //                                            .dir_TX
		output wire        tx_qsys_conduit_drv_en_TX,                                 //                                            .drv_en_TX
		output wire        tr_qsys_conduit_drv_en_TR,                                 //                             tr_qsys_conduit.drv_en_TR
		output wire        tr_qsys_conduit_dir_TR,                                    //                                            .dir_TR
		output wire        tr_qsys_conduit_counter_en_TR,                             //                                            .counter_en_TR
		output wire [15:0] tr_qsys_conduit_period_TR,                                 //                                            .period_TR
		input  wire        tr_qsys_conduit_dir_AUTO,                                  //                                            .dir_AUTO
		input  wire        tr_qsys_conduit_dir_MANUAL,                                //                                            .dir_MANUAL
		input  wire        tr_qsys_conduit_auto,                                      //                                            .auto
		input  wire        tr_qsys_conduit_enable_AUTO,                               //                                            .enable_AUTO
		input  wire        tr_qsys_conduit_enable_MANUAL,                             //                                            .enable_MANUAL
		input  wire [15:0] tr_qsys_conduit_period_AUTO,                               //                                            .period_AUTO
		input  wire        tr_qsys_conduit_count_MANUAL,                              //                                            .count_MANUAL
		input  wire [15:0] tr_qsys_conduit_period_MANUAL,                             //                                            .period_MANUAL
		output wire        tr_auto_qsys_conduit_enable_AUTO,                          //                        tr_auto_qsys_conduit.enable_AUTO
		output wire        tr_auto_qsys_conduit_dir_AUTO,                             //                                            .dir_AUTO
		output wire [31:0] tr_auto_qsys_conduit_period_AUTO,                          //                                            .period_AUTO
		input  wire        tr_auto_qsys_conduit_data_valid_TR,                        //                                            .data_valid_TR
		input  wire        tr_auto_qsys_conduit_tr_mode,                              //                                            .tr_mode
		input  wire [11:0] tr_auto_qsys_conduit_x_set,                                //                                            .x_set
		input  wire [15:0] tr_auto_qsys_conduit_x,                                    //                                            .x
		input  wire [15:0] tr_auto_qsys_conduit_dx1,                                  //                                            .dx1
		input  wire [15:0] tr_auto_qsys_conduit_dx2,                                  //                                            .dx2
		input  wire [15:0] tr_auto_qsys_conduit_F1,                                   //                                            .F1
		input  wire [15:0] tr_auto_qsys_conduit_F2,                                   //                                            .F2
		input  wire [15:0] tr_auto_qsys_conduit_DZ_TR,                                //                                            .DZ_TR
		input  wire [19:0] tr_auto_qsys_conduit_k_TR,                                 //                                            .k_TR
		input  wire [15:0] tr_auto_qsys_conduit_L,                                    //                                            .L
		input  wire [31:0] tr_manual_qsys_conduit_count_N,                            //                      tr_manual_qsys_conduit.count_N
		input  wire [31:0] tr_manual_qsys_conduit_PULSE_NUMBER,                       //                                            .PULSE_NUMBER
		output wire        tr_manual_qsys_conduit_enable_MANUAL,                      //                                            .enable_MANUAL
		input  wire        tr_manual_qsys_conduit_stop,                               //                                            .stop
		input  wire        tr_manual_qsys_conduit_start_N,                            //                                            .start_N
		input  wire        tr_manual_qsys_conduit_start                               //                                            .start
	);

	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [15:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_debugaccess;                               // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;             // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire  [31:0] mm_interconnect_0_pio_led_s1_writedata;                    // mm_interconnect_0:pio_led_s1_writedata -> pio_led:writedata
	wire   [1:0] mm_interconnect_0_pio_led_s1_address;                      // mm_interconnect_0:pio_led_s1_address -> pio_led:address
	wire         mm_interconnect_0_pio_led_s1_chipselect;                   // mm_interconnect_0:pio_led_s1_chipselect -> pio_led:chipselect
	wire         mm_interconnect_0_pio_led_s1_write;                        // mm_interconnect_0:pio_led_s1_write -> pio_led:write_n
	wire  [31:0] mm_interconnect_0_pio_led_s1_readdata;                     // pio_led:readdata -> mm_interconnect_0:pio_led_s1_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [15:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;             // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire  [12:0] mm_interconnect_0_onchip_memory2_s1_address;               // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;            // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                 // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         mm_interconnect_0_onchip_memory2_s1_write;                 // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;              // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;            // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;       // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;         // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;           // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;             // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;              // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;          // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] cpu_d_irq_irq;                                             // irq_mapper:sender_irq -> cpu:d_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [cpu:reset_n, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, mux_qsys_0:rst, onchip_memory2:reset, pio_led:reset_n, pulse_qsys_0:rst, rst_translator:in_reset, sysid:reset_n, tp_qsys_0:rst, tr_auto_qsys_0:rst, tr_manual_qsys_0:rst, tr_qsys_0:rst, tx_qsys_0:rst]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu:reset_req, onchip_memory2:reset_req, rst_translator:reset_req_in]
	wire         cpu_jtag_debug_module_reset_reset;                         // cpu:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> commands_parameters_qsys_0:rst

	master_cpu cpu (
		.clk                                   (clk_50),                                              //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	master_jtag_uart jtag_uart (
		.clk            (clk_50),                                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	master_onchip_memory2 onchip_memory2 (
		.clk        (clk_50),                                         //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)              //       .reset_req
	);

	master_pio_led pio_led (
		.clk        (clk_50),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_s1_readdata),   //                    .readdata
		.out_port   (pio_led_external_connection_export)       // external_connection.export
	);

	master_sysid sysid (
		.clock    (clk_50),                                         //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	COMMANDS_PARAMETERS #(
		.WIDTH_C_P (16)
	) commands_parameters_qsys_0 (
		.clk              (clk_50),                                                    //            clock.clk
		.avs_s0_address   (commands_parameters_qsys_0_s0_address),                     //               s0.address
		.avs_s0_writedata (commands_parameters_qsys_0_s0_writedata),                   //                 .writedata
		.avs_s0_readdata  (commands_parameters_qsys_0_s0_readdata),                    //                 .readdata
		.avs_s0_write     (commands_parameters_qsys_0_s0_write),                       //                 .write
		.avs_s0_read      (commands_parameters_qsys_0_s0_read),                        //                 .read
		.rst              (rst_controller_001_reset_out_reset),                        //            reset.reset
		.start            (commands_parameters_qsys_0_conduit_comm_par_start),         // conduit_comm_par.export
		.start_N          (commands_parameters_qsys_0_conduit_comm_par_start_N),       //                 .export
		.auto             (commands_parameters_qsys_0_conduit_comm_par_auto),          //                 .export
		.stop             (commands_parameters_qsys_0_conduit_comm_par_stop),          //                 .export
		.fi_phm           (commands_parameters_qsys_0_conduit_comm_par_fi_phm),        //                 .export
		.detuning         (commands_parameters_qsys_0_conduit_comm_par_detuning),      //                 .export
		.syncpulse        (commands_parameters_qsys_0_conduit_comm_par_syncpulse),     //                 .export
		.TURN_ON_RF       (commands_parameters_qsys_0_conduit_comm_par_TURN_ON_RF),    //                 .export
		.d_fi_gate2       (commands_parameters_qsys_0_conduit_comm_par_d_fi_gate2),    //                 .export
		.d_i_gate2        (commands_parameters_qsys_0_conduit_comm_par_d_i_gate2),     //                 .export
		.dx2              (commands_parameters_qsys_0_conduit_comm_par_dx2),           //                 .export
		.dx1              (commands_parameters_qsys_0_conduit_comm_par_dx1),           //                 .export
		.DZ_TP            (commands_parameters_qsys_0_conduit_comm_par_DZ_TP),         //                 .export
		.DZ_TX            (commands_parameters_qsys_0_conduit_comm_par_DZ_TX),         //                 .export
		.PULSE_NUMBER     (commands_parameters_qsys_0_conduit_comm_par_PULSE_NUMBER),  //                 .export
		.DZ_TR            (commands_parameters_qsys_0_conduit_comm_par_DZ_TR),         //                 .export
		.period_MANUAL    (commands_parameters_qsys_0_conduit_comm_par_period_MANUAL), //                 .export
		.L                (commands_parameters_qsys_0_conduit_comm_par_L),             //                 .export
		.F2               (commands_parameters_qsys_0_conduit_comm_par_F2),            //                 .export
		.F1               (commands_parameters_qsys_0_conduit_comm_par_F1),            //                 .export
		.count_MANUAL     (commands_parameters_qsys_0_conduit_comm_par_count_MANUAL),  //                 .export
		.dir_MANUAL       (commands_parameters_qsys_0_conduit_comm_par_dir_MANUAL),    //                 .export
		.tp               (commands_parameters_qsys_0_conduit_comm_par_tp),            //                 .export
		.tx               (commands_parameters_qsys_0_conduit_comm_par_tx),            //                 .export
		.tr               (commands_parameters_qsys_0_conduit_comm_par_tr)             //                 .export
	);

	TR_MANUAL #(
		.WIDTH_MANUAL (16)
	) tr_manual_qsys_0 (
		.clk           (clk_50),                               //             clock.clk
		.rst           (rst_controller_reset_out_reset),       //             reset.reset
		.count_N       (tr_manual_qsys_conduit_count_N),       // conduit_tr_manual.export
		.PULSE_NUMBER  (tr_manual_qsys_conduit_PULSE_NUMBER),  //                  .export
		.enable_MANUAL (tr_manual_qsys_conduit_enable_MANUAL), //                  .export
		.stop          (tr_manual_qsys_conduit_stop),          //                  .export
		.start_N       (tr_manual_qsys_conduit_start_N),       //                  .export
		.start         (tr_manual_qsys_conduit_start)          //                  .export
	);

	TR_AUTO #(
		.WIDTH_IN   (12),
		.WIDTH_AUTO (16)
	) tr_auto_qsys_0 (
		.clk           (clk_50),                             //           clock.clk
		.rst           (rst_controller_reset_out_reset),     //           reset.reset
		.enable_AUTO   (tr_auto_qsys_conduit_enable_AUTO),   // conduit_tr_auto.export
		.dir_AUTO      (tr_auto_qsys_conduit_dir_AUTO),      //                .export
		.period_AUTO   (tr_auto_qsys_conduit_period_AUTO),   //                .export
		.data_valid_TR (tr_auto_qsys_conduit_data_valid_TR), //                .export
		.tr_mode       (tr_auto_qsys_conduit_tr_mode),       //                .export
		.x_set         (tr_auto_qsys_conduit_x_set),         //                .export
		.x             (tr_auto_qsys_conduit_x),             //                .export
		.dx1           (tr_auto_qsys_conduit_dx1),           //                .export
		.dx2           (tr_auto_qsys_conduit_dx2),           //                .export
		.F1            (tr_auto_qsys_conduit_F1),            //                .export
		.F2            (tr_auto_qsys_conduit_F2),            //                .export
		.DZ_TR         (tr_auto_qsys_conduit_DZ_TR),         //                .export
		.k_TR          (tr_auto_qsys_conduit_k_TR),          //                .export
		.L             (tr_auto_qsys_conduit_L)              //                .export
	);

	TR #(
		.WIDTH_TR (16)
	) tr_qsys_0 (
		.clk           (clk_50),                         //      clock.clk
		.rst           (rst_controller_reset_out_reset), //      reset.reset
		.drv_en_TR     (tr_qsys_conduit_drv_en_TR),      // conduit_tr.export
		.dir_TR        (tr_qsys_conduit_dir_TR),         //           .export
		.counter_en_TR (tr_qsys_conduit_counter_en_TR),  //           .export
		.period_TR     (tr_qsys_conduit_period_TR),      //           .export
		.dir_AUTO      (tr_qsys_conduit_dir_AUTO),       //           .export
		.dir_MANUAL    (tr_qsys_conduit_dir_MANUAL),     //           .export
		.auto          (tr_qsys_conduit_auto),           //           .export
		.enable_AUTO   (tr_qsys_conduit_enable_AUTO),    //           .export
		.enable_MANUAL (tr_qsys_conduit_enable_MANUAL),  //           .export
		.period_AUTO   (tr_qsys_conduit_period_AUTO),    //           .export
		.count_MANUAL  (tr_qsys_conduit_count_MANUAL),   //           .export
		.period_MANUAL (tr_qsys_conduit_period_MANUAL)   //           .export
	);

	TX #(
		.WIDTH_TX (16)
	) tx_qsys_0 (
		.clk           (clk_50),                         //      clock.clk
		.rst           (rst_controller_reset_out_reset), //      reset.reset
		.syncpulse     (tx_qsys_conduit_syncpulse),      // conduit_tx.export
		.k_TX          (tx_qsys_conduit_k_TX),           //           .export
		.d_i_gate2     (tx_qsys_conduit_d_i_gate2),      //           .export
		.DZ_TX         (tx_qsys_conduit_DZ_TX),          //           .export
		.L             (tx_qsys_conduit_L),              //           .export
		.F2            (tx_qsys_conduit_F2),             //           .export
		.F1            (tx_qsys_conduit_F1),             //           .export
		.i_fid_TX      (tx_qsys_conduit_i_fid_TX),       //           .export
		.i_set         (tx_qsys_conduit_i_set),          //           .export
		.tx_mode       (tx_qsys_conduit_tx_mode),        //           .export
		.i_fid         (tx_qsys_conduit_i_fid),          //           .export
		.data_valid_TX (tx_qsys_conduit_data_valid_TX),  //           .export
		.period_TX     (tx_qsys_conduit_period_TX),      //           .export
		.dir_TX        (tx_qsys_conduit_dir_TX),         //           .export
		.drv_en_TX     (tx_qsys_conduit_drv_en_TX)       //           .export
	);

	TP #(
		.WIDTH_TP (16)
	) tp_qsys_0 (
		.rst           (rst_controller_reset_out_reset), //      reset.reset
		.k_TP          (tp_qsys_conduit_k_TP),           // conduit_tp.export
		.d_fi_gate2    (tp_qsys_conduit_d_fi_gate2),     //           .export
		.L             (tp_qsys_conduit_L),              //           .export
		.DZ_TP         (tp_qsys_conduit_DZ_TP),          //           .export
		.F2            (tp_qsys_conduit_F2),             //           .export
		.F1            (tp_qsys_conduit_F1),             //           .export
		.detuning      (tp_qsys_conduit_detuning),       //           .export
		.fi_set        (tp_qsys_conduit_fi_set),         //           .export
		.fi_phm        (tp_qsys_conduit_fi_phm),         //           .export
		.tp_mode       (tp_qsys_conduit_tp_mode),        //           .export
		.data_valid_TP (tp_qsys_conduit_data_valid_TP),  //           .export
		.period_TP     (tp_qsys_conduit_period_TP),      //           .export
		.dir_TP        (tp_qsys_conduit_dir_TP),         //           .export
		.drv_en_TP     (tp_qsys_conduit_drv_en_TP),      //           .export
		.clk           (clk_50)                          //      clock.clk
	);

	MUX #(
		.WIDTH_MUX (16)
	) mux_qsys_0 (
		.clk           (clk_50),                         //       clock.clk
		.rst           (rst_controller_reset_out_reset), //       reset.reset
		.drv_period    (mux_qsys_conduit_drv_period),    // conduit_mux.export
		.drv_dir       (mux_qsys_conduit_drv_dir),       //            .export
		.enable        (mux_qsys_conduit_enable),        //            .export
		.counter_en    (mux_qsys_conduit_counter_en),    //            .export
		.period_TR     (mux_qsys_conduit_period_TR),     //            .export
		.period_TX     (mux_qsys_conduit_period_TX),     //            .export
		.period_TP     (mux_qsys_conduit_period_TP),     //            .export
		.detuning      (mux_qsys_conduit_detuning),      //            .export
		.fi_phm        (mux_qsys_conduit_fi_phm),        //            .export
		.tr            (mux_qsys_conduit_tr),            //            .export
		.tx            (mux_qsys_conduit_tx),            //            .export
		.tp            (mux_qsys_conduit_tp),            //            .export
		.dir_TX        (mux_qsys_conduit_dir_TX),        //            .export
		.dir_TR        (mux_qsys_conduit_dir_TR),        //            .export
		.dir_TP        (mux_qsys_conduit_dir_TP),        //            .export
		.drv_en_TR     (mux_qsys_conduit_drv_en_TR),     //            .export
		.drv_en_TX     (mux_qsys_conduit_drv_en_TX),     //            .export
		.drv_en_TP     (mux_qsys_conduit_drv_en_TP),     //            .export
		.counter_en_TR (mux_qsys_conduit_counter_en_TR), //            .export
		.syncpulse     (mux_qsys_conduit_syncpulse)      //            .export
	);

	PULSE #(
		.WIDTH (16)
	) pulse_qsys_0 (
		.clk          (clk_50),                          //         clock.clk
		.rst          (rst_controller_reset_out_reset),  //         reset.reset
		.drv_pulse    (pulse_qsys_conduit_drv_pulse),    // conduit_pulse.export
		.drv_dir      (pulse_qsys_conduit_drv_dir),      //              .export
		.enable       (pulse_qsys_conduit_enable),       //              .export
		.counter_en   (pulse_qsys_conduit_counter_en),   //              .export
		.drv_period   (pulse_qsys_conduit_drv_period),   //              .export
		.PULSE_NUMBER (pulse_qsys_conduit_PULSE_NUMBER)  //              .export
	);

	master_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                          (clk_50),                                                    //                        clk_50_clk.clk
		.cpu_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // cpu_reset_n_reset_bridge_in_reset.reset
		.cpu_data_master_address                 (cpu_data_master_address),                                   //                   cpu_data_master.address
		.cpu_data_master_waitrequest             (cpu_data_master_waitrequest),                               //                                  .waitrequest
		.cpu_data_master_byteenable              (cpu_data_master_byteenable),                                //                                  .byteenable
		.cpu_data_master_read                    (cpu_data_master_read),                                      //                                  .read
		.cpu_data_master_readdata                (cpu_data_master_readdata),                                  //                                  .readdata
		.cpu_data_master_write                   (cpu_data_master_write),                                     //                                  .write
		.cpu_data_master_writedata               (cpu_data_master_writedata),                                 //                                  .writedata
		.cpu_data_master_debugaccess             (cpu_data_master_debugaccess),                               //                                  .debugaccess
		.cpu_instruction_master_address          (cpu_instruction_master_address),                            //            cpu_instruction_master.address
		.cpu_instruction_master_waitrequest      (cpu_instruction_master_waitrequest),                        //                                  .waitrequest
		.cpu_instruction_master_read             (cpu_instruction_master_read),                               //                                  .read
		.cpu_instruction_master_readdata         (cpu_instruction_master_readdata),                           //                                  .readdata
		.cpu_jtag_debug_module_address           (mm_interconnect_0_cpu_jtag_debug_module_address),           //             cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write             (mm_interconnect_0_cpu_jtag_debug_module_write),             //                                  .write
		.cpu_jtag_debug_module_read              (mm_interconnect_0_cpu_jtag_debug_module_read),              //                                  .read
		.cpu_jtag_debug_module_readdata          (mm_interconnect_0_cpu_jtag_debug_module_readdata),          //                                  .readdata
		.cpu_jtag_debug_module_writedata         (mm_interconnect_0_cpu_jtag_debug_module_writedata),         //                                  .writedata
		.cpu_jtag_debug_module_byteenable        (mm_interconnect_0_cpu_jtag_debug_module_byteenable),        //                                  .byteenable
		.cpu_jtag_debug_module_waitrequest       (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),       //                                  .waitrequest
		.cpu_jtag_debug_module_debugaccess       (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),       //                                  .debugaccess
		.jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //       jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                  .write
		.jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                  .read
		.jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                  .readdata
		.jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                  .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                  .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                  .chipselect
		.onchip_memory2_s1_address               (mm_interconnect_0_onchip_memory2_s1_address),               //                 onchip_memory2_s1.address
		.onchip_memory2_s1_write                 (mm_interconnect_0_onchip_memory2_s1_write),                 //                                  .write
		.onchip_memory2_s1_readdata              (mm_interconnect_0_onchip_memory2_s1_readdata),              //                                  .readdata
		.onchip_memory2_s1_writedata             (mm_interconnect_0_onchip_memory2_s1_writedata),             //                                  .writedata
		.onchip_memory2_s1_byteenable            (mm_interconnect_0_onchip_memory2_s1_byteenable),            //                                  .byteenable
		.onchip_memory2_s1_chipselect            (mm_interconnect_0_onchip_memory2_s1_chipselect),            //                                  .chipselect
		.onchip_memory2_s1_clken                 (mm_interconnect_0_onchip_memory2_s1_clken),                 //                                  .clken
		.pio_led_s1_address                      (mm_interconnect_0_pio_led_s1_address),                      //                        pio_led_s1.address
		.pio_led_s1_write                        (mm_interconnect_0_pio_led_s1_write),                        //                                  .write
		.pio_led_s1_readdata                     (mm_interconnect_0_pio_led_s1_readdata),                     //                                  .readdata
		.pio_led_s1_writedata                    (mm_interconnect_0_pio_led_s1_writedata),                    //                                  .writedata
		.pio_led_s1_chipselect                   (mm_interconnect_0_pio_led_s1_chipselect),                   //                                  .chipselect
		.sysid_control_slave_address             (mm_interconnect_0_sysid_control_slave_address),             //               sysid_control_slave.address
		.sysid_control_slave_readdata            (mm_interconnect_0_sysid_control_slave_readdata)             //                                  .readdata
	);

	master_irq_mapper irq_mapper (
		.clk           (clk_50),                         //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (clk_50),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.clk            (clk_50),                             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
