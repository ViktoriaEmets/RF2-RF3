module MASTER  // совсем не то написано 
(
	input                           clk,
	output wire			start,
   output wire			stop,
   output wire			start_N,
                
	output wire			avto,
	output wire			drv_pulse,
	output wire			drv_dir
	
);

endmodule 
