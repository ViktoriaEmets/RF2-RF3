`timescale 10ns/10ns
module Test();
 
reg          clk_50MHz,
             rst,
             data_valid,
        	    syncpulse,
        	    tr_mode,
        	    tx_mode,
        	    tp_mode; 
        	    
integer      i_set = 50,
             i_fid_TX = 100,
        	    d_i_gate2 = 95,
             DZ_TX = 25,
             
        	    fi_set = 70,
        	    d_fi_gate2 = 65,
        	    DZ_TP = 25,
        	    detuning = 70;
        	    
        	      
        	    
integer      L = 16,
             x_set = 35,
             DZ_TR  = 100,
        	    dx1 = 150,
        	    dx2 = 400,
        	    F1 = 6000,
        	    F2 = 50000;

wire [31:0]  L_conn,
             F1_conn,
             F2_conn;   	    
        	    
//--------------------------------- CLK -------------------------------------------------------------------------
initial
begin
  clk_50MHz = 0;
  forever
  clk_50MHz = #10!clk_50MHz;
end
//--------------------------------------------------------------------------------------------------------------


//----------------------- RST -----------------------------------------------------------------------------------
initial
begin
  rst =0;
  #5100 rst=1;
  #3000 rst=0;
end
//---------------------------------------------------------------------------------------------------------------


//------------------------------ DATA_VALID ----------------------------------------------------------------------
initial
begin
  data_valid=0;
 forever
  begin
      data_valid=0;
    repeat(4)
    @(posedge clk_50MHz);
      data_valid=1;
    @(posedge clk_50MHz);
  end
end
//---------------------------------------------------------------------------------------------------------------


//------------------------------------------- DELAY ------------------------------------------------------------
task delay;
input integer T;
repeat (T)
@(posedge clk_50MHz);
endtask
//-------------------------------------------------------------------------------------------------------------


//---------------------------------------- syncpulse -----------------------------------------------------------
initial
begin
  syncpulse =0;
  #170000 syncpulse=1;
  #10 syncpulse=0;
end
//----------------------------------------------------------------------------------------------------------------


//------------------------------ find k -----------------------------------------------------------------------------
integer k_TR;
initial
begin
  k_TR=((F2 - F1)/(dx2 - dx1)) * L;
  $display("k_TR = %d", k_TR);
end  
//-----------------------------------------------
integer k_TX;
initial
begin
  k_TX=((F2 - F1)/(d_i_gate2 - DZ_TX)) * L;
  $display("k_TX = %d", k_TX);
end  
//------------------------------------------------
integer k_TP;
initial
begin
  k_TP=((F2 - F1)/(d_fi_gate2 - DZ_TP)) * L;
  $display("k_TP = %d", k_TP);
end        	    
//--------------------------------------------------------------------------------------------------------------- 


//-------------------------- tr_mode ------------------------------------------------------------------------------------
initial
begin
  tr_mode = 0;
  #30000 tr_mode = 1;
  #50000 tr_mode = 0;
  #20000 tr_mode = 1;
end
//--------------------------- tx_mode ------------------------
initial
begin
  tx_mode = 0;
  #170000 tx_mode = 1;
  #500000 tx_mode = 0;
  #200000 tx_mode = 1;
end
//--------------------------- tp_mode --------------------------
initial
begin
  tp_mode = 0;
  #220000 tp_mode = 1;
  #500000 tp_mode = 0;
  #200000 tp_mode = 1;
end
//--------------------------------------------------------------------------------------------------------------------------


//----------------------------------- X --------------------------------------------------------------------------------
parameter    F=450;
reg [15:0]   x;
always @(posedge data_valid)
begin
        if (tr_mode == 0)
          begin
            x = 500;
          end 
   
        else 
          begin
            if (x > 0)
   	           begin 
                    x = x - 1;
               end
 	          else 
                begin 
                  while(x < F)
                    x = x + 1;
                end
            end
    end
//--------------------------------------------------------------------------------------------------------------------------


//----------------------------------- i_fid --------------------------------------------------------------------------------
reg [15:0]   i_fid;
always @(posedge clk_50MHz)
begin
  if(syncpulse || tx_mode == 1)
    begin  
      if (i_fid <= 7000)
        begin
          i_fid <= i_fid + 1; 
        end  
      else
        begin
          i_fid <=i_fid;
        end  
    end
  else
    begin
     i_fid <= 10; 
    end
end      
//--------------------------------------------------------------------------------------------------------------------------


//----------------------------------- fi_phm --------------------------------------------------------------------------------
reg [15:0]   fi_phm;
always @(posedge clk_50MHz)
begin
        if (tp_mode == 0)
          begin
            fi_phm = 180;
          end 
   
        else 
          begin
            if (fi_phm > 0)
   	           begin 
                    fi_phm = fi_phm - 1;
               end
 	          else 
                begin 
                    fi_phm = 0;
                end
            end
    end
//--------------------------------------------------------------------------------------------------------------------------

//--------------------------------------------------------------------------------------------------------------------------
TR TR_Test
(
  .clk                (clk_50MHz),
  .data_valid         (data_valid), 
  .tr_mode            (tr_mode), 
  .rst                (rst), 

  .x                  (x), 
  .x_set              (x_set),
  .dx1                (dx1), 
  .dx2                (dx2),
  .DZ_TR              (DZ_TR),
  .L                  (L_conn),
  .F2                 (F2),
  .F1                 (F1),
  .k_TR               (k_TR) 
);

TX TX_Test
(
  .clk                (clk_50MHz), 
  .tx_mode            (tx_mode), 
  .rst                (rst), 

  .i_fid              (i_fid),          
  .i_set              (i_set),           
  .i_fid_TX           (i_fid_TX),
  .syncpulse          (syncpulse),
  .DZ_TX              (DZ_TX),
  .d_i_gate2          (d_i_gate2),
  
  .L                  (L_conn),
  .F2                 (F2_conn),
  .F1                 (F1_conn) 
);

TP TP_Test
(
  .clk                (clk_50MHz), 
  .tp_mode            (tp_mode), 
  .rst                (rst), 
  
  .fi_phm             (fi_phm),
  .fi_set             (fi_set),
  .detuning           (detuning),
  .DZ_TP              (DZ_TP),
  .d_fi_gate2         (d_fi_gate2),
  
  .L                  (L_conn),
  .F2                 (F2_conn),
  .F1                 (F1_conn)  
);

PULSE PULSE_test
(
  .clk                (clk_50MHz),  
  .rst                (rst), 
  .drv_pulse          (drv_pulse)
);


endmodule
